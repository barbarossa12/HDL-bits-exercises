// https://hdlbits.01xz.net/wiki/Adder100
module top_module( 
    input [99:0] a, b,
    input cin,
    output cout,
    output [99:0] sum );

    wire [100:0] result;
    assign result = {1'b0, a} + {1'b0, b} + cin;
    assign sum = result[99:0];
    assign cout = result[100];
endmodule


// a simpler solution would be to do the following
// assign {cout, sum} = a + b + cin;
//
